module baud_gen (
    input clk,
    input [16:0] baud_gen
);

    